package spi_package;

   `include "spi_transaction.sv"
   `include "spi_generator.sv"
   `include "spi_driver.sv"
   `include "spi_monitor.sv"
   `include "spi_scoreboard.sv"
   `include "spi_environment.sv"

endpackage